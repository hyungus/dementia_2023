
module gameover (clk, reset, gameend);

input clk, reset, gameend;


wire clk, reset, gameend;
